module clk_dic()
  int
  reg
  wire
  
